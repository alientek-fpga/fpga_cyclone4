library verilog;
use verilog.vl_types.all;
entity sdram_tb is
end sdram_tb;
