library verilog;
use verilog.vl_types.all;
entity sdr is
    generic(
        tCK             : real    := 6.000000;
        tCK3_min        : real    := 6.000000;
        tCK2_min        : real    := 10.000000;
        tCK1_min        : real    := 20.000000;
        tAC3            : real    := 5.400000;
        tAC2            : real    := 7.500000;
        tAC1            : real    := 17.000000;
        tHZ3            : real    := 5.400000;
        tHZ2            : real    := 7.500000;
        tHZ1            : real    := 17.000000;
        tOH             : real    := 3.000000;
        tMRD            : real    := 2.000000;
        tRAS            : real    := 42.000000;
        tRC             : real    := 60.000000;
        tRFC            : real    := 60.000000;
        tRCD            : real    := 18.000000;
        tRP             : real    := 18.000000;
        tRRD            : real    := 2.000000;
        tWRa            : real    := 6.000000;
        tWRm            : real    := 12.000000;
        ADDR_BITS       : integer := 12;
        ROW_BITS        : integer := 12;
        COL_BITS        : integer := 9;
        DQ_BITS         : integer := 16;
        DM_BITS         : integer := 2;
        BA_BITS         : integer := 2;
        mem_sizes       : vl_notype
    );
    port(
        Dq              : inout  vl_logic_vector;
        Addr            : in     vl_logic_vector;
        Ba              : in     vl_logic_vector;
        Clk             : in     vl_logic;
        Cke             : in     vl_logic;
        Cs_n            : in     vl_logic;
        Ras_n           : in     vl_logic;
        Cas_n           : in     vl_logic;
        We_n            : in     vl_logic;
        Dqm             : in     vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of tCK : constant is 1;
    attribute mti_svvh_generic_type of tCK3_min : constant is 1;
    attribute mti_svvh_generic_type of tCK2_min : constant is 1;
    attribute mti_svvh_generic_type of tCK1_min : constant is 1;
    attribute mti_svvh_generic_type of tAC3 : constant is 1;
    attribute mti_svvh_generic_type of tAC2 : constant is 1;
    attribute mti_svvh_generic_type of tAC1 : constant is 1;
    attribute mti_svvh_generic_type of tHZ3 : constant is 1;
    attribute mti_svvh_generic_type of tHZ2 : constant is 1;
    attribute mti_svvh_generic_type of tHZ1 : constant is 1;
    attribute mti_svvh_generic_type of tOH : constant is 1;
    attribute mti_svvh_generic_type of tMRD : constant is 1;
    attribute mti_svvh_generic_type of tRAS : constant is 1;
    attribute mti_svvh_generic_type of tRC : constant is 1;
    attribute mti_svvh_generic_type of tRFC : constant is 1;
    attribute mti_svvh_generic_type of tRCD : constant is 1;
    attribute mti_svvh_generic_type of tRP : constant is 1;
    attribute mti_svvh_generic_type of tRRD : constant is 1;
    attribute mti_svvh_generic_type of tWRa : constant is 1;
    attribute mti_svvh_generic_type of tWRm : constant is 1;
    attribute mti_svvh_generic_type of ADDR_BITS : constant is 1;
    attribute mti_svvh_generic_type of ROW_BITS : constant is 1;
    attribute mti_svvh_generic_type of COL_BITS : constant is 1;
    attribute mti_svvh_generic_type of DQ_BITS : constant is 1;
    attribute mti_svvh_generic_type of DM_BITS : constant is 1;
    attribute mti_svvh_generic_type of BA_BITS : constant is 1;
    attribute mti_svvh_generic_type of mem_sizes : constant is 3;
end sdr;
