//****************************************Copyright (c)***********************************//
//����֧�֣�www.openedv.com
//�Ա����̣�http://openedv.taobao.com 
//��ע΢�Ź���ƽ̨΢�źţ�"����ԭ��"����ѻ�ȡFPGA & STM32���ϡ�
//��Ȩ���У�����ؾ���
//Copyright(C) ����ԭ�� 2018-2028
//All rights reserved	                               
//----------------------------------------------------------------------------------------
// File name:          tb_top_key_beep
// Last modified Date:  2018��5��7��14:33:28
// Last Version:        V1.1
// Descriptions:        ��������
//----------------------------------------------------------------------------------------
// Created by:          ����ԭ��
// Created date:        2018��5��7��14:33:33
// Version:             V1.0
// Descriptions:        The original version
//
//----------------------------------------------------------------------------------------
// Modified by:		    ����ԭ��
// Modified date:	    2018/4/24 9:56:36
// Version:			    V1.1
// Descriptions:	    �������Ʒ���������ģ��
//
//----------------------------------------------------------------------------------------
//****************************************************************************************//
`timescale 1 ns/ 1 ns
module tb_top_key_beep();

//parameter define
parameter T = 20;

//reg define
reg  key;
reg  sys_clk;
reg  sys_rst_n;
reg  key_value;

// wire define                                               
wire beep;

//*****************************************************
//**                    main code                  
//*****************************************************

//���źų�ʼֵ
initial begin
    key                          <= 1'b1;
    sys_clk                      <= 1'b0;
    sys_rst_n                    <= 1'b0; 
    #20           sys_rst_n      <= 1'b1;  //�ڵ�20ns��ʱ��λ�ź��ź����� 
    #30           key            <= 1'b0;  //�ڵ�50ns��ʱ���°���
    #20           key            <= 1'b1;  //ģ�ⶶ��
    #20           key            <= 1'b0;  //ģ�ⶶ��
    #20           key            <= 1'b1;  //ģ�ⶶ��
    #20           key            <= 1'b0;  //ģ�ⶶ��
    #170          key            <= 1'b1;  //�ڵ�300ns��ʱ���ɿ�����
    #20           key            <= 1'b0;  //ģ�ⶶ��
    #20           key            <= 1'b1;  //ģ�ⶶ��
    #20           key            <= 1'b0;  //ģ�ⶶ��
    #20           key            <= 1'b1;  //ģ�ⶶ��
    #170          key            <= 1'b0;  //�ڵ�550ns��ʱ���ٴΰ��°���
    #20           key            <= 1'b1;  //ģ�ⶶ��
    #20           key            <= 1'b0;  //ģ�ⶶ��
    #20           key            <= 1'b1;  //ģ�ⶶ��
    #20           key            <= 1'b0;  //ģ�ⶶ��
    #170          key            <= 1'b1;  //�ڵ�800ns��ʱ���ɿ�����
    #20           key            <= 1'b0;  //ģ�ⶶ��
    #20           key            <= 1'b1;  //ģ�ⶶ��
    #20           key            <= 1'b0;  //ģ�ⶶ��
    #20           key            <= 1'b1;  //ģ�ⶶ��
end

//50Mhz��ʱ�ӣ�������Ϊ1/50Mhz=20ns,����ÿ10ns����ƽȡ��һ��  
 always # (T/2) sys_clk <= ~sys_clk;

//����key_beepģ��                        
top_key_beep u1 (
	.beep(beep),
	.key(key),
	.sys_clk(sys_clk),
	.sys_rst_n(sys_rst_n)
);           
                                       
endmodule
