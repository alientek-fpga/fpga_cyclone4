//****************************************Copyright (c)***********************************//
//技术支持：www.openedv.com
//淘宝店铺：http://openedv.taobao.com 
//关注微信公众平台微信号："正点原子"，免费获取FPGA & STM32资料。
//版权所有，盗版必究。
//Copyright(C) 正点原子 2018-2028
//All rights reserved	                               
//----------------------------------------------------------------------------------------
// File name:           lcd_display
// Last modified Date:  2018/1/30 11:12:36
// Last Version:        V1.1
// Descriptions:        RGB LCD字符显示模块
//----------------------------------------------------------------------------------------
// Created by:          正点原子
// Created date:        2018/1/29 10:55:56
// Version:             V1.0
// Descriptions:        The original version
//
//----------------------------------------------------------------------------------------
// Modified by:		    正点原子
// Modified date:	    2018/1/30 11:12:36
// Version:			    V1.1
// Descriptions:	    在RGB LCD上显示汉字”正点原子”
//
//----------------------------------------------------------------------------------------
//****************************************************************************************//

module lcd_display(
    input             lcd_clk,                  //lcd驱动时钟
    input             sys_rst_n,                //复位信号
    
    input      [10:0] pixel_xpos,               //像素点横坐标
    input      [10:0] pixel_ypos,               //像素点纵坐标    
    output reg [15:0] pixel_data                //像素点数据,
    );    

//parameter define    
parameter  H_DISP = 11'd800;                    //分辨率——行
parameter  V_DISP = 11'd480;                    //分辨率——列

localparam POS_X  = 11'd336;                    //字符区域起始点横坐标
localparam POS_Y  = 11'd224;                    //字符区域起始点纵坐标
localparam WIDTH  = 11'd128;                    //字符区域宽度
localparam HEIGHT = 11'd32;                     //字符区域高度
localparam RED    = 16'b11111_000000_00000;     //屏幕背景色
localparam BLUE   = 16'b00000_000000_11111;     //字符颜色
localparam BLACK  = 16'b00000_000000_00000;     //字符区域背景色

//reg define
reg  [127:0] char[31:0];                        //字符数组

//wire define   
wire [10:0] x_cnt;
wire [10:0] y_cnt;

//*****************************************************
//**                    main code
//*****************************************************
assign x_cnt = pixel_xpos - POS_X;              //像素点相对于字符区域起始点水平坐标
assign y_cnt = pixel_ypos - POS_Y;              //像素点相对于字符区域起始点竖直坐标

//给字符数组赋值，显示汉字“正点原子”，汉字大小为32*32
always @(posedge lcd_clk) begin
    char[0 ]  <= 128'h00000000000000000000000000000000;
    char[1 ]  <= 128'h00000000000000000000000000000000;
    char[2 ]  <= 128'h00000000000100000000002000000000;
    char[3 ]  <= 128'h000000380001800002000070000000C0;
    char[4 ]  <= 128'h0000007C0001800003FFFFF803FFFFE0;
    char[5 ]  <= 128'h0FFFFFFE0001800003006000000001E0;
    char[6 ]  <= 128'h0001E000000180600300600000000300;
    char[7 ]  <= 128'h0001E0000001FFF00300C00000000600;
    char[8 ]  <= 128'h0001E000000180000310804000001800;
    char[9 ]  <= 128'h0001E00000018000031FFFE000003000;
    char[10]  <= 128'h0001E00000018000031800400001C000;
    char[11]  <= 128'h0181E00000018000031800400001C000;
    char[12]  <= 128'h01E1E000018181800318004000018000;
    char[13]  <= 128'h01F1E00001FFFFC0031FFFC000018010;
    char[14]  <= 128'h01E1E0E0018001800318004000018038;
    char[15]  <= 128'h01E1FFF001800180031800403FFFFFFC;
    char[16]  <= 128'h01E1E018018001800318004000018000;
    char[17]  <= 128'h01E1E000018001800218004000018000;
    char[18]  <= 128'h01E1E00001800180021FFFC000018000;
    char[19]  <= 128'h01E1E000018001800210304000018000;
    char[20]  <= 128'h01E1E00001FFFF800200300000018000;
    char[21]  <= 128'h01E1E000018001800606300000018000;
    char[22]  <= 128'h01E1E000018001000607370000018000;
    char[23]  <= 128'h01E1E00000000000060E31C000018000;
    char[24]  <= 128'h01E1E000001000400418307000018000;
    char[25]  <= 128'h01E1E000020830600430303800018000;
    char[26]  <= 128'h01E1E038020C18300860301800018000;
    char[27]  <= 128'h01E1E07C060E18180883700800018000;
    char[28]  <= 128'h7FFFFFFE0C0618181100F008003F8000;
    char[29]  <= 128'h000000001C0408182000600000070000;
    char[30]  <= 128'h00000000000000000000000000020000;
    char[31]  <= 128'h00000000000000000000000000000000;
end

//给不同的区域绘制不同的颜色
always @(posedge lcd_clk or negedge sys_rst_n) begin         
    if (!sys_rst_n) 
        pixel_data <= BLACK;
    else begin
        if((pixel_xpos >= POS_X) && (pixel_xpos < POS_X + WIDTH)
          && (pixel_ypos >= POS_Y) && (pixel_ypos < POS_Y + HEIGHT)) begin
            if(char[y_cnt][11'd127 - x_cnt])
                pixel_data <= BLUE;             //绘制字符为蓝色
            else
                pixel_data <= BLACK;            //绘制字符区域背景为黑色      
        end
        else
            pixel_data <= RED;                  //绘制屏幕背景为红色
    end
end

endmodule 